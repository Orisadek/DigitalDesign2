//
// Verilog Module Lab2AlonOri_lib.matmul
//
// Created:
//          by - orisad.UNKNOWN (TOMER)
//          at - 19:03:27 02/15/2024
//
// using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
//

`resetall
`timescale 1ns/10ps
module matmul(clk_i,rst_ni,psel_i,penable_i,pwrite_i,pstrb_i,pwdata_i,paddr_i,pready_o,pslverr_o,prdata_o,busy_o);





endmodule
